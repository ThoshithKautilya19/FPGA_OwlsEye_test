`timescale 1 ns / 1 ps

module AESL_deadlock_report_unit #( parameter PROC_NUM = 4 ) (
    input reset,
    input clock,
    input [PROC_NUM - 1:0] dl_in_vec,
    output dl_detect_out,
    output reg [PROC_NUM - 1:0] origin,
    output token_clear);
   
    // FSM states
    localparam ST_IDLE = 2'b0;
    localparam ST_DL_DETECTED = 2'b1;
    localparam ST_DL_REPORT = 2'b10;

    reg [1:0] CS_fsm;
    reg [1:0] NS_fsm;
    reg [PROC_NUM - 1:0] dl_detect_reg;
    reg [PROC_NUM - 1:0] dl_done_reg;
    reg [PROC_NUM - 1:0] origin_reg;
    reg [PROC_NUM - 1:0] dl_in_vec_reg;
    integer i;
    integer fp;

    // FSM State machine
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            CS_fsm <= ST_IDLE;
        end
        else begin
            CS_fsm <= NS_fsm;
        end
    end
    always @ (CS_fsm or dl_in_vec or dl_detect_reg or dl_done_reg or dl_in_vec or origin_reg) begin
        NS_fsm = CS_fsm;
        case (CS_fsm)
            ST_IDLE : begin
                if (|dl_in_vec) begin
                    NS_fsm = ST_DL_DETECTED;
                end
            end
            ST_DL_DETECTED: begin
                // has unreported deadlock cycle
                if (dl_detect_reg != dl_done_reg) begin
                    NS_fsm = ST_DL_REPORT;
                end
            end
            ST_DL_REPORT: begin
                if (|(dl_in_vec & origin_reg)) begin
                    NS_fsm = ST_DL_DETECTED;
                end
            end
        endcase
    end

    // dl_detect_reg record the procs that first detect deadlock
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            dl_detect_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_IDLE) begin
                dl_detect_reg <= dl_in_vec;
            end
        end
    end

    // dl_detect_out keeps in high after deadlock detected
    assign dl_detect_out = |dl_detect_reg;

    // dl_done_reg record the cycles has been reported
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            dl_done_reg <= 'b0;
        end
        else begin
            if ((CS_fsm == ST_DL_REPORT) && (|(dl_in_vec & dl_detect_reg) == 'b1)) begin
                dl_done_reg <= dl_done_reg | dl_in_vec;
            end
        end
    end

    // clear token once a cycle is done
    assign token_clear = (CS_fsm == ST_DL_REPORT) ? ((|(dl_in_vec & origin_reg)) ? 'b1 : 'b0) : 'b0;

    // origin_reg record the current cycle start id
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            origin_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                origin_reg <= origin;
            end
        end
    end
   
    // origin will be valid for only one cycle
    always @ (CS_fsm or dl_detect_reg or dl_done_reg) begin
        origin = 'b0;
        if (CS_fsm == ST_DL_DETECTED) begin
            for (i = 0; i < PROC_NUM; i = i + 1) begin
                if (dl_detect_reg[i] & ~dl_done_reg[i] & ~(|origin)) begin
                    origin = 'b1 << i;
                end
            end
        end
    end
    
    // dl_in_vec_reg record the current cycle dl_in_vec
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            dl_in_vec_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                dl_in_vec_reg <= origin;
            end
            else if (CS_fsm == ST_DL_REPORT) begin
                dl_in_vec_reg <= dl_in_vec;
            end
        end
    end
    
    // get the first valid proc index in dl vector
    function integer proc_index(input [PROC_NUM - 1:0] dl_vec);
        begin
            proc_index = 0;
            for (i = 0; i < PROC_NUM; i = i + 1) begin
                if (dl_vec[i]) begin
                    proc_index = i;
                end
            end
        end
    endfunction

    // get the proc path based on dl vector
    function [1128:0] proc_path(input [PROC_NUM - 1:0] dl_vec);
        integer index;
        begin
            index = proc_index(dl_vec);
            case (index)
                0 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.mem_read36130_U0";
                end
                1 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0";
                end
                2 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0";
                end
                3 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_line_U0";
                end
                4 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0";
                end
                5 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0";
                end
                6 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0";
                end
                7 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0";
                end
                8 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0";
                end
                9 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0";
                end
                10 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0";
                end
                11 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0";
                end
                12 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1";
                end
                13 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1";
                end
                14 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0";
                end
                15 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0";
                end
                16 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2";
                end
                17 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2";
                end
                18 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0";
                end
                19 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0";
                end
                20 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3";
                end
                21 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3";
                end
                22 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_glue_U0";
                end
                23 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias199_U0";
                end
                24 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias200_U0";
                end
                25 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias201_U0";
                end
                26 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias202_U0";
                end
                27 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0";
                end
                28 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_in_U0";
                end
                29 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0";
                end
                30 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0";
                end
                31 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu203_U0";
                end
                32 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu204_U0";
                end
                33 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu205_U0";
                end
                34 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu206_U0";
                end
                35 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu207_U0";
                end
                36 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu208_U0";
                end
                37 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu209_U0";
                end
                38 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu210_U0";
                end
                39 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu211_U0";
                end
                40 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu212_U0";
                end
                41 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu213_U0";
                end
                42 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu214_U0";
                end
                43 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu215_U0";
                end
                44 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu216_U0";
                end
                45 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu217_U0";
                end
                46 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu218_U0";
                end
                47 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0";
                end
                48 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0";
                end
                49 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0";
                end
                50 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.mem_write_U0";
                end
                51 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_reload_weights_fu_524.mem_read_U0";
                end
                52 : begin
                    proc_path = "fpgaconvnet_ip.Block_proc_U0.grp_reload_weights_fu_524.weights_reloading_U0";
                end
                default : begin
                    proc_path = "unknown";
                end
            endcase
        end
    endfunction

    // print the headlines of deadlock detection
    task print_dl_head;
        begin
            $display("\n//////////////////////////////////////////////////////////////////////////////");
            $display("// ERROR!!! DEADLOCK DETECTED at %0t ns! SIMULATION WILL BE STOPPED! //", $time);
            $display("//////////////////////////////////////////////////////////////////////////////");
            fp = $fopen("deadlock_db.dat", "w");
        end
    endtask

    // print the start of a cycle
    task print_cycle_start(input reg [1128:0] proc_path, input integer cycle_id);
        begin
            $display("/////////////////////////");
            $display("// Dependence cycle %0d:", cycle_id);
            $display("// (1): Process: %0s", proc_path);
            $fdisplay(fp, "Dependence_Cycle_ID %0d", cycle_id);
            $fdisplay(fp, "Dependence_Process_ID 1");
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print the end of deadlock detection
    task print_dl_end(input integer num);
        begin
            $display("////////////////////////////////////////////////////////////////////////");
            $display("// Totally %0d cycles detected!", num);
            $display("////////////////////////////////////////////////////////////////////////");
            $fdisplay(fp, "Dependence_Cycle_Number %0d", num);
            $fclose(fp);
        end
    endtask

    // print one proc component in the cycle
    task print_cycle_proc_comp(input reg [1128:0] proc_path, input integer cycle_comp_id);
        begin
            $display("// (%0d): Process: %0s", cycle_comp_id, proc_path);
            $fdisplay(fp, "Dependence_Process_ID %0d", cycle_comp_id);
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print one channel component in the cycle
    task print_cycle_chan_comp(input [PROC_NUM - 1:0] dl_vec1, input [PROC_NUM - 1:0] dl_vec2);
        reg [1096:0] chan_path;
        integer index1;
        integer index2;
        begin
            index1 = proc_index(dl_vec1);
            index2 = proc_index(dl_vec2);
            case (index1)
                0 : begin
                    case(index2)
                    2: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.mem_read36130_U0.in_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.in_0_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.in_0_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.in_0_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    50: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.mem_read36130_U0.weights_reloading_in_3_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.weights_reloading_in_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.weights_reloading_in_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.weights_reloading_in_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.mem_read36130_U0.out_hw_V_offset_out_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_hw_V_offset_c_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_hw_V_offset_c_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_hw_V_offset_c_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.start_for_mem_wriFfa_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.mem_write_U0.ap_done)) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.start_for_mem_wriFfa_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.mem_write_U0.ap_done)) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    1: begin
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.start_for_Conv_0_U0_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.ap_done)) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.start_for_Conv_0_U0_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.ap_done)) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    endcase
                end
                1 : begin
                    case(index2)
                    0: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_line_U0.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.in_0_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.in_0_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.in_0_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.start_for_Conv_0_U0_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.ap_idle))) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.start_for_Conv_0_U0_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.ap_idle))) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    28: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias199_U0.grp_bias_fu_28.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias200_U0.grp_bias372_fu_28.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias201_U0.grp_bias371_fu_28.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias202_U0.grp_bias370_fu_28.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    27: begin
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.start_for_Conv_0_Gfk_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.ap_done)) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.start_for_Conv_0_Gfk_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.ap_done)) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    endcase
                end
                2 : begin
                    case(index2)
                    0: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_line_U0.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.in_0_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.in_0_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.in_0_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    5: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.out_V_V1_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.out_V_V2_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.out_V_V3_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.out_V_V4_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.out_V_V25_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.out_V_V255_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.out_V_V256_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.out_V_V257_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.out_V_V258_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.out_V_V26_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.out_V_V269_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.out_V_V2610_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.out_V_V2611_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.out_V_V2612_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.out_V_V27_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.out_V_V2713_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.out_V_V2714_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.out_V_V2715_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.out_V_V2716_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.out_V_V28_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.out_V_V2817_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.out_V_V2818_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.out_V_V2819_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.out_V_V2820_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_qcK_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.ap_done)) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_qcK_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.ap_done)) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    endcase
                end
                3 : begin
                    case(index2)
                    4: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_line_U0.frame_buffer_0_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_line_U0.frame_buffer_0_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_line_U0.frame_buffer_0_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_line_U0.frame_buffer_0_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_line_U0.frame_buffer_0_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_line_U0.frame_buffer_1_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_line_U0.frame_buffer_1_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_line_U0.frame_buffer_1_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_line_U0.frame_buffer_1_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_line_U0.frame_buffer_1_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_line_U0.frame_buffer_2_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_line_U0.frame_buffer_2_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_line_U0.frame_buffer_2_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_line_U0.frame_buffer_2_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_line_U0.frame_buffer_2_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_line_U0.frame_buffer_3_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_line_U0.frame_buffer_3_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_line_U0.frame_buffer_3_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_line_U0.frame_buffer_3_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_line_U0.frame_buffer_3_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_line_U0.frame_buffer_4_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_line_U0.frame_buffer_4_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_line_U0.frame_buffer_4_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_line_U0.frame_buffer_4_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_line_U0.frame_buffer_4_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.start_for_slidingcud_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.ap_done)) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.start_for_slidingcud_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.ap_done)) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    endcase
                end
                4 : begin
                    case(index2)
                    3: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.frame_buffer_0_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.frame_buffer_0_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.frame_buffer_0_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.frame_buffer_0_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.frame_buffer_0_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_0_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.frame_buffer_1_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.frame_buffer_1_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.frame_buffer_1_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.frame_buffer_1_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.frame_buffer_1_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_1_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.frame_buffer_2_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.frame_buffer_2_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.frame_buffer_2_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.frame_buffer_2_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.frame_buffer_2_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_2_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.frame_buffer_3_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.frame_buffer_3_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.frame_buffer_3_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.frame_buffer_3_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.frame_buffer_3_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_3_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.frame_buffer_4_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.frame_buffer_4_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.frame_buffer_4_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.frame_buffer_4_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.frame_buffer_4_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.frame_buffer_4_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.start_for_slidingcud_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.ap_idle))) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.start_for_slidingcud_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_sliding_windo_U0.grp_sliding_window_fu_66.sliding_window_out_U0.ap_idle))) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    endcase
                end
                5 : begin
                    case(index2)
                    2: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.in_V_V1_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.in_V_V2_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.in_V_V3_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.in_V_V4_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_0_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.in_V_V15_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.in_V_V16_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.in_V_V17_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.in_V_V18_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.in_V_V19_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_1_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.in_V_V210_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.in_V_V211_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.in_V_V212_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.in_V_V213_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.in_V_V214_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_2_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.in_V_V315_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.in_V_V316_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.in_V_V317_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.in_V_V318_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.in_V_V319_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_3_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.in_V_V420_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.in_V_V421_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.in_V_V422_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.in_V_V423_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.in_V_V424_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.sw_out_0_4_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_qcK_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.ap_idle))) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_qcK_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.ap_idle))) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    6: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_0_0_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_0_0_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_0_0_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_0_0_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_0_0_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_0_1_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_0_1_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_0_1_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_0_1_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_0_1_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_0_2_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_0_2_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_0_2_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_0_2_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_0_2_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_0_3_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_0_3_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_0_3_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_0_3_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_0_3_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_0_4_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_0_4_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_0_4_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_0_4_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_0_4_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_rcU_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.ap_done)) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_rcU_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.ap_done)) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    10: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_1_0_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_1_0_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_1_0_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_1_0_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_1_0_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_1_1_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_1_1_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_1_1_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_1_1_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_1_1_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_1_2_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_1_2_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_1_2_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_1_2_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_1_2_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_1_3_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_1_3_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_1_3_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_1_3_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_1_3_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_1_4_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_1_4_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_1_4_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_1_4_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_1_4_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_sc4_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.ap_done)) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_sc4_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.ap_done)) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    14: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_2_0_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_2_0_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_2_0_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_2_0_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_2_0_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_2_1_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_2_1_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_2_1_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_2_1_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_2_1_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_2_2_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_2_2_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_2_2_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_2_2_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_2_2_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_2_3_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_2_3_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_2_3_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_2_3_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_2_3_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_2_4_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_2_4_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_2_4_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_2_4_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_2_4_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_tde_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.ap_done)) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_tde_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.ap_done)) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    18: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_3_0_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_3_0_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_3_0_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_3_0_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_3_0_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_3_1_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_3_1_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_3_1_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_3_1_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_3_1_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_3_2_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_3_2_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_3_2_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_3_2_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_3_2_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_3_3_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_3_3_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_3_3_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_3_3_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_3_3_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_3_4_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_3_4_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_3_4_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_3_4_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_fork194_U0.grp_fork_r_fu_264.out_3_4_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_udo_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.ap_done)) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_udo_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.ap_done)) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    endcase
                end
                6 : begin
                    case(index2)
                    5: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.in_V_V1_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.in_V_V2_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.in_V_V3_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.in_V_V4_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_0_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.in_V_V15_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.in_V_V16_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.in_V_V17_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.in_V_V18_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.in_V_V19_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_1_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.in_V_V210_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.in_V_V211_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.in_V_V212_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.in_V_V213_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.in_V_V214_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_2_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.in_V_V315_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.in_V_V316_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.in_V_V317_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.in_V_V318_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.in_V_V319_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_3_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.in_V_V420_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.in_V_V421_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.in_V_V422_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.in_V_V423_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.in_V_V424_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_0_4_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_rcU_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.ap_idle))) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_rcU_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.ap_idle))) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    22: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.conv_out_0_0_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.conv_out_0_0_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.conv_out_0_0_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_vdy_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_glue_U0.ap_done)) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_vdy_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_glue_U0.ap_done)) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    endcase
                end
                7 : begin
                    case(index2)
                    8: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.window_stream_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.window_stream_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.window_stream_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.window_stream_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.window_stream_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.window_stream_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.window_stream_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.window_stream_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.window_stream_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_8_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_8_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_8_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.window_stream_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_9_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_9_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_9_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.window_stream_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_10_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_10_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_10_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.window_stream_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_11_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_11_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_11_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.window_stream_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_12_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_12_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_12_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.window_stream_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_13_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_13_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_13_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.window_stream_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_14_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_14_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_14_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.window_stream_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_15_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_15_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_15_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.window_stream_16_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_16_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_16_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_16_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.window_stream_17_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.window_stream_18_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.window_stream_19_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.window_stream_20_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.window_stream_21_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.window_stream_22_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.window_stream_23_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.window_stream_24_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.weight_stream_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.weight_stream_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.weight_stream_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.weight_stream_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.weight_stream_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.weight_stream_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.weight_stream_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.weight_stream_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.weight_stream_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_8_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_8_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_8_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.weight_stream_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_9_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_9_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_9_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.weight_stream_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_10_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_10_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_10_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.weight_stream_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_11_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_11_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_11_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.weight_stream_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_12_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_12_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_12_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.weight_stream_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_13_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_13_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_13_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.weight_stream_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_14_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_14_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_14_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.weight_stream_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_15_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_15_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_15_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.weight_stream_16_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_16_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_16_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_16_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.weight_stream_17_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.weight_stream_18_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.weight_stream_19_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.weight_stream_20_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.weight_stream_21_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.weight_stream_22_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.weight_stream_23_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_intr_U0.weight_stream_24_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.start_for_conv_mueOg_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.ap_done)) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.start_for_conv_mueOg_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.ap_done)) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    endcase
                end
                8 : begin
                    case(index2)
                    7: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.window_stream_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.window_stream_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.window_stream_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.window_stream_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.window_stream_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.window_stream_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.window_stream_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.window_stream_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.window_stream_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_8_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_8_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_8_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.window_stream_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_9_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_9_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_9_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.window_stream_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_10_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_10_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_10_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.window_stream_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_11_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_11_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_11_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.window_stream_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_12_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_12_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_12_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.window_stream_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_13_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_13_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_13_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.window_stream_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_14_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_14_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_14_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.window_stream_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_15_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_15_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_15_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.window_stream_16_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_16_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_16_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_16_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.window_stream_17_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.window_stream_18_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.window_stream_19_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.window_stream_20_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.window_stream_21_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.window_stream_22_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.window_stream_23_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.window_stream_24_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.weight_stream_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.weight_stream_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.weight_stream_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.weight_stream_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.weight_stream_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.weight_stream_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.weight_stream_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.weight_stream_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.weight_stream_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_8_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_8_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_8_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.weight_stream_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_9_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_9_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_9_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.weight_stream_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_10_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_10_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_10_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.weight_stream_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_11_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_11_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_11_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.weight_stream_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_12_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_12_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_12_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.weight_stream_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_13_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_13_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_13_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.weight_stream_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_14_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_14_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_14_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.weight_stream_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_15_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_15_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_15_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.weight_stream_16_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_16_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_16_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_16_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.weight_stream_17_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.weight_stream_18_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.weight_stream_19_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.weight_stream_20_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.weight_stream_21_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.weight_stream_22_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.weight_stream_23_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.weight_stream_24_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.start_for_conv_mueOg_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.ap_idle))) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.start_for_conv_mueOg_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.ap_idle))) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    9: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.acc_stream_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.acc_stream_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.acc_stream_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.acc_stream_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.acc_stream_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.acc_stream_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.acc_stream_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.acc_stream_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.acc_stream_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_8_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_8_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_8_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.acc_stream_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_9_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_9_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_9_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.acc_stream_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_10_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_10_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_10_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.acc_stream_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_11_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_11_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_11_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.acc_stream_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_12_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_12_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_12_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.acc_stream_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_13_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_13_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_13_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.acc_stream_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_14_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_14_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_14_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.acc_stream_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_15_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_15_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_15_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.acc_stream_16_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_16_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_16_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_16_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.acc_stream_17_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.acc_stream_18_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.acc_stream_19_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.acc_stream_20_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.acc_stream_21_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.acc_stream_22_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.acc_stream_23_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_mul_U0.acc_stream_24_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.start_for_conv_acfYi_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.ap_done)) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.start_for_conv_acfYi_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.ap_done)) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    endcase
                end
                9 : begin
                    case(index2)
                    8: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.acc_stream_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.acc_stream_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.acc_stream_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.acc_stream_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.acc_stream_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.acc_stream_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.acc_stream_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.acc_stream_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.acc_stream_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_8_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_8_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_8_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.acc_stream_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_9_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_9_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_9_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.acc_stream_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_10_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_10_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_10_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.acc_stream_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_11_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_11_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_11_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.acc_stream_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_12_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_12_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_12_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.acc_stream_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_13_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_13_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_13_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.acc_stream_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_14_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_14_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_14_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.acc_stream_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_15_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_15_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_15_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.acc_stream_16_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_16_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_16_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_16_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.acc_stream_17_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.acc_stream_18_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.acc_stream_19_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.acc_stream_20_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.acc_stream_21_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.acc_stream_22_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.acc_stream_23_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.acc_stream_24_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.start_for_conv_acfYi_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.ap_idle))) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.start_for_conv_acfYi_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.conv_acc_U0.ap_idle))) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    endcase
                end
                10 : begin
                    case(index2)
                    5: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.in_V_V1_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.in_V_V2_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.in_V_V3_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.in_V_V4_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_0_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.in_V_V15_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.in_V_V16_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.in_V_V17_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.in_V_V18_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.in_V_V19_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_1_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.in_V_V210_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.in_V_V211_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.in_V_V212_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.in_V_V213_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.in_V_V214_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_2_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.in_V_V315_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.in_V_V316_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.in_V_V317_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.in_V_V318_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.in_V_V319_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_3_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.in_V_V420_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.in_V_V421_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.in_V_V422_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.in_V_V423_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.in_V_V424_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_1_4_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_sc4_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.ap_idle))) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_sc4_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.ap_idle))) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    22: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.conv_out_0_1_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.conv_out_0_1_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.conv_out_0_1_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                11 : begin
                    case(index2)
                    12: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.window_stream_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.window_stream_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.window_stream_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.window_stream_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.window_stream_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.window_stream_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.window_stream_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.window_stream_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.window_stream_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_8_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_8_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_8_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.window_stream_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_9_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_9_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_9_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.window_stream_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_10_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_10_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_10_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.window_stream_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_11_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_11_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_11_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.window_stream_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_12_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_12_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_12_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.window_stream_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_13_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_13_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_13_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.window_stream_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_14_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_14_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_14_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.window_stream_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_15_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_15_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_15_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.window_stream_16_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_16_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_16_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_16_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.window_stream_17_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.window_stream_18_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.window_stream_19_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.window_stream_20_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.window_stream_21_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.window_stream_22_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.window_stream_23_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.window_stream_24_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.window_stream_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.weight_stream_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.weight_stream_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.weight_stream_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.weight_stream_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.weight_stream_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.weight_stream_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.weight_stream_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.weight_stream_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.weight_stream_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_8_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_8_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_8_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.weight_stream_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_9_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_9_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_9_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.weight_stream_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_10_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_10_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_10_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.weight_stream_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_11_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_11_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_11_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.weight_stream_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_12_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_12_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_12_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.weight_stream_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_13_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_13_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_13_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.weight_stream_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_14_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_14_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_14_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.weight_stream_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_15_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_15_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_15_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.weight_stream_16_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_16_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_16_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_16_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.weight_stream_17_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.weight_stream_18_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.weight_stream_19_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.weight_stream_20_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.weight_stream_21_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.weight_stream_22_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.weight_stream_23_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_intr369_U0.weight_stream_24_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.weight_stream_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.start_for_conv_mug8j_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.ap_done)) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.start_for_conv_mug8j_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.ap_done)) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    endcase
                end
                12 : begin
                    case(index2)
                    7: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.window_stream_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.window_stream_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.window_stream_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.window_stream_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.window_stream_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.window_stream_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.window_stream_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.window_stream_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.window_stream_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_8_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_8_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_8_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.window_stream_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_9_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_9_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_9_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.window_stream_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_10_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_10_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_10_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.window_stream_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_11_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_11_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_11_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.window_stream_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_12_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_12_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_12_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.window_stream_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_13_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_13_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_13_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.window_stream_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_14_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_14_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_14_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.window_stream_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_15_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_15_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_15_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.window_stream_16_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_16_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_16_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_16_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.window_stream_17_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.window_stream_18_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.window_stream_19_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.window_stream_20_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.window_stream_21_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.window_stream_22_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.window_stream_23_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.window_stream_24_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.weight_stream_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.weight_stream_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.weight_stream_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.weight_stream_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.weight_stream_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.weight_stream_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.weight_stream_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.weight_stream_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.weight_stream_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_8_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_8_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_8_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.weight_stream_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_9_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_9_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_9_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.weight_stream_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_10_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_10_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_10_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.weight_stream_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_11_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_11_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_11_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.weight_stream_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_12_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_12_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_12_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.weight_stream_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_13_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_13_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_13_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.weight_stream_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_14_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_14_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_14_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.weight_stream_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_15_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_15_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_15_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.weight_stream_16_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_16_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_16_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_16_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.weight_stream_17_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.weight_stream_18_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.weight_stream_19_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.weight_stream_20_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.weight_stream_21_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.weight_stream_22_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.weight_stream_23_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.weight_stream_24_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    9: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.acc_stream_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.acc_stream_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.acc_stream_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.acc_stream_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.acc_stream_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.acc_stream_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.acc_stream_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.acc_stream_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.acc_stream_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_8_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_8_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_8_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.acc_stream_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_9_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_9_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_9_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.acc_stream_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_10_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_10_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_10_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.acc_stream_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_11_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_11_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_11_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.acc_stream_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_12_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_12_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_12_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.acc_stream_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_13_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_13_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_13_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.acc_stream_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_14_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_14_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_14_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.acc_stream_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_15_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_15_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_15_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.acc_stream_16_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_16_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_16_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_16_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.acc_stream_17_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.acc_stream_18_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.acc_stream_19_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.acc_stream_20_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.acc_stream_21_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.acc_stream_22_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.acc_stream_23_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.acc_stream_24_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    11: begin
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.start_for_conv_mug8j_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.ap_idle))) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.start_for_conv_mug8j_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_mul_U1_1.ap_idle))) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    13: begin
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.start_for_conv_achbi_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.ap_done)) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.start_for_conv_achbi_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.ap_done)) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    endcase
                end
                13 : begin
                    case(index2)
                    8: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.acc_stream_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.acc_stream_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.acc_stream_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.acc_stream_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.acc_stream_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.acc_stream_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.acc_stream_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.acc_stream_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.acc_stream_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_8_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_8_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_8_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.acc_stream_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_9_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_9_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_9_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.acc_stream_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_10_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_10_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_10_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.acc_stream_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_11_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_11_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_11_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.acc_stream_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_12_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_12_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_12_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.acc_stream_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_13_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_13_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_13_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.acc_stream_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_14_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_14_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_14_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.acc_stream_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_15_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_15_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_15_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.acc_stream_16_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_16_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_16_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_16_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.acc_stream_17_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.acc_stream_18_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.acc_stream_19_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.acc_stream_20_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.acc_stream_21_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.acc_stream_22_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.acc_stream_23_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.acc_stream_24_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    12: begin
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.start_for_conv_achbi_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.ap_idle))) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.start_for_conv_achbi_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv196_U0.grp_conv368_fu_126.conv_acc_U1_1.ap_idle))) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    endcase
                end
                14 : begin
                    case(index2)
                    5: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.in_V_V1_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.in_V_V2_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.in_V_V3_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.in_V_V4_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_0_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.in_V_V15_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.in_V_V16_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.in_V_V17_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.in_V_V18_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.in_V_V19_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_1_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.in_V_V210_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.in_V_V211_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.in_V_V212_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.in_V_V213_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.in_V_V214_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_2_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.in_V_V315_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.in_V_V316_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.in_V_V317_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.in_V_V318_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.in_V_V319_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_3_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.in_V_V420_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.in_V_V421_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.in_V_V422_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.in_V_V423_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.in_V_V424_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_2_4_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_tde_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.ap_idle))) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_tde_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.ap_idle))) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    22: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.conv_out_0_2_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.conv_out_0_2_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.conv_out_0_2_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                15 : begin
                    case(index2)
                    16: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.window_stream_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.window_stream_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.window_stream_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.window_stream_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.window_stream_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.window_stream_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.window_stream_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.window_stream_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.window_stream_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_8_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_8_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_8_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.window_stream_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_9_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_9_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_9_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.window_stream_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_10_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_10_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_10_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.window_stream_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_11_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_11_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_11_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.window_stream_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_12_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_12_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_12_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.window_stream_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_13_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_13_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_13_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.window_stream_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_14_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_14_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_14_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.window_stream_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_15_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_15_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_15_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.window_stream_16_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_16_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_16_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_16_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.window_stream_17_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.window_stream_18_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.window_stream_19_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.window_stream_20_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.window_stream_21_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.window_stream_22_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.window_stream_23_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.window_stream_24_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.window_stream_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.weight_stream_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.weight_stream_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.weight_stream_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.weight_stream_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.weight_stream_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.weight_stream_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.weight_stream_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.weight_stream_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.weight_stream_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_8_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_8_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_8_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.weight_stream_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_9_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_9_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_9_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.weight_stream_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_10_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_10_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_10_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.weight_stream_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_11_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_11_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_11_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.weight_stream_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_12_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_12_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_12_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.weight_stream_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_13_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_13_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_13_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.weight_stream_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_14_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_14_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_14_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.weight_stream_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_15_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_15_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_15_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.weight_stream_16_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_16_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_16_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_16_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.weight_stream_17_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.weight_stream_18_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.weight_stream_19_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.weight_stream_20_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.weight_stream_21_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.weight_stream_22_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.weight_stream_23_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_intr367_U0.weight_stream_24_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.weight_stream_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.start_for_conv_muibs_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.ap_done)) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.start_for_conv_muibs_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.ap_done)) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    endcase
                end
                16 : begin
                    case(index2)
                    7: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.window_stream_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.window_stream_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.window_stream_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.window_stream_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.window_stream_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.window_stream_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.window_stream_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.window_stream_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.window_stream_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_8_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_8_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_8_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.window_stream_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_9_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_9_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_9_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.window_stream_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_10_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_10_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_10_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.window_stream_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_11_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_11_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_11_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.window_stream_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_12_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_12_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_12_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.window_stream_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_13_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_13_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_13_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.window_stream_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_14_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_14_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_14_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.window_stream_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_15_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_15_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_15_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.window_stream_16_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_16_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_16_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_16_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.window_stream_17_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.window_stream_18_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.window_stream_19_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.window_stream_20_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.window_stream_21_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.window_stream_22_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.window_stream_23_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.window_stream_24_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.weight_stream_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.weight_stream_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.weight_stream_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.weight_stream_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.weight_stream_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.weight_stream_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.weight_stream_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.weight_stream_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.weight_stream_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_8_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_8_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_8_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.weight_stream_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_9_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_9_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_9_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.weight_stream_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_10_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_10_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_10_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.weight_stream_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_11_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_11_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_11_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.weight_stream_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_12_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_12_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_12_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.weight_stream_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_13_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_13_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_13_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.weight_stream_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_14_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_14_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_14_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.weight_stream_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_15_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_15_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_15_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.weight_stream_16_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_16_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_16_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_16_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.weight_stream_17_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.weight_stream_18_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.weight_stream_19_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.weight_stream_20_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.weight_stream_21_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.weight_stream_22_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.weight_stream_23_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.weight_stream_24_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    9: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.acc_stream_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.acc_stream_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.acc_stream_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.acc_stream_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.acc_stream_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.acc_stream_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.acc_stream_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.acc_stream_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.acc_stream_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_8_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_8_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_8_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.acc_stream_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_9_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_9_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_9_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.acc_stream_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_10_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_10_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_10_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.acc_stream_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_11_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_11_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_11_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.acc_stream_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_12_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_12_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_12_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.acc_stream_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_13_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_13_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_13_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.acc_stream_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_14_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_14_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_14_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.acc_stream_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_15_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_15_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_15_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.acc_stream_16_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_16_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_16_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_16_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.acc_stream_17_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.acc_stream_18_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.acc_stream_19_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.acc_stream_20_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.acc_stream_21_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.acc_stream_22_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.acc_stream_23_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.acc_stream_24_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    15: begin
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.start_for_conv_muibs_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.ap_idle))) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.start_for_conv_muibs_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_mul_U2_2.ap_idle))) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    17: begin
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.start_for_conv_acjbC_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.ap_done)) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.start_for_conv_acjbC_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.ap_done)) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    endcase
                end
                17 : begin
                    case(index2)
                    8: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.acc_stream_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.acc_stream_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.acc_stream_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.acc_stream_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.acc_stream_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.acc_stream_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.acc_stream_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.acc_stream_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.acc_stream_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_8_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_8_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_8_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.acc_stream_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_9_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_9_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_9_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.acc_stream_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_10_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_10_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_10_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.acc_stream_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_11_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_11_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_11_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.acc_stream_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_12_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_12_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_12_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.acc_stream_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_13_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_13_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_13_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.acc_stream_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_14_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_14_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_14_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.acc_stream_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_15_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_15_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_15_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.acc_stream_16_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_16_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_16_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_16_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.acc_stream_17_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.acc_stream_18_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.acc_stream_19_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.acc_stream_20_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.acc_stream_21_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.acc_stream_22_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.acc_stream_23_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.acc_stream_24_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    16: begin
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.start_for_conv_acjbC_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.ap_idle))) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.start_for_conv_acjbC_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv197_U0.grp_conv366_fu_126.conv_acc_U2_2.ap_idle))) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    endcase
                end
                18 : begin
                    case(index2)
                    5: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.in_V_V1_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.in_V_V2_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.in_V_V3_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.in_V_V4_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_0_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.in_V_V15_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.in_V_V16_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.in_V_V17_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.in_V_V18_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.in_V_V19_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_1_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.in_V_V210_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.in_V_V211_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.in_V_V212_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.in_V_V213_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.in_V_V214_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_2_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.in_V_V315_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.in_V_V316_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.in_V_V317_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.in_V_V318_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.in_V_V319_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_3_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.in_V_V420_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.in_V_V421_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.in_V_V422_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.in_V_V423_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.in_V_V424_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.fork_out_0_3_4_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_udo_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.ap_idle))) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_udo_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.ap_idle))) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    22: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.conv_out_0_3_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.conv_out_0_3_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.conv_out_0_3_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                19 : begin
                    case(index2)
                    20: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.window_stream_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.window_stream_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.window_stream_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.window_stream_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.window_stream_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.window_stream_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.window_stream_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.window_stream_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.window_stream_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_8_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_8_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_8_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.window_stream_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_9_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_9_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_9_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.window_stream_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_10_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_10_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_10_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.window_stream_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_11_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_11_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_11_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.window_stream_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_12_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_12_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_12_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.window_stream_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_13_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_13_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_13_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.window_stream_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_14_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_14_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_14_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.window_stream_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_15_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_15_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_15_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.window_stream_16_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_16_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_16_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_16_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.window_stream_17_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.window_stream_18_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.window_stream_19_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.window_stream_20_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.window_stream_21_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.window_stream_22_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.window_stream_23_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.window_stream_24_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.window_stream_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.weight_stream_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.weight_stream_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.weight_stream_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.weight_stream_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.weight_stream_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.weight_stream_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.weight_stream_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.weight_stream_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.weight_stream_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_8_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_8_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_8_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.weight_stream_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_9_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_9_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_9_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.weight_stream_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_10_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_10_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_10_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.weight_stream_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_11_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_11_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_11_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.weight_stream_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_12_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_12_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_12_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.weight_stream_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_13_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_13_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_13_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.weight_stream_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_14_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_14_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_14_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.weight_stream_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_15_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_15_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_15_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.weight_stream_16_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_16_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_16_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_16_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.weight_stream_17_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.weight_stream_18_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.weight_stream_19_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.weight_stream_20_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.weight_stream_21_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.weight_stream_22_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.weight_stream_23_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_intr365_U0.weight_stream_24_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.weight_stream_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.start_for_conv_mukbM_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.ap_done)) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.start_for_conv_mukbM_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.ap_done)) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    endcase
                end
                20 : begin
                    case(index2)
                    7: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.window_stream_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.window_stream_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.window_stream_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.window_stream_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.window_stream_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.window_stream_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.window_stream_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.window_stream_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.window_stream_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_8_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_8_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_8_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.window_stream_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_9_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_9_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_9_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.window_stream_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_10_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_10_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_10_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.window_stream_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_11_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_11_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_11_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.window_stream_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_12_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_12_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_12_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.window_stream_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_13_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_13_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_13_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.window_stream_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_14_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_14_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_14_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.window_stream_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_15_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_15_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_15_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.window_stream_16_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_16_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_16_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_16_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.window_stream_17_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.window_stream_18_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.window_stream_19_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.window_stream_20_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.window_stream_21_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.window_stream_22_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.window_stream_23_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.window_stream_24_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.window_stream_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.weight_stream_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.weight_stream_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.weight_stream_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.weight_stream_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.weight_stream_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.weight_stream_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.weight_stream_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.weight_stream_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.weight_stream_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_8_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_8_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_8_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.weight_stream_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_9_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_9_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_9_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.weight_stream_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_10_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_10_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_10_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.weight_stream_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_11_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_11_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_11_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.weight_stream_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_12_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_12_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_12_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.weight_stream_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_13_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_13_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_13_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.weight_stream_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_14_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_14_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_14_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.weight_stream_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_15_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_15_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_15_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.weight_stream_16_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_16_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_16_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_16_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.weight_stream_17_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.weight_stream_18_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.weight_stream_19_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.weight_stream_20_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.weight_stream_21_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.weight_stream_22_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.weight_stream_23_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.weight_stream_24_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.weight_stream_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    9: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.acc_stream_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.acc_stream_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.acc_stream_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.acc_stream_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.acc_stream_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.acc_stream_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.acc_stream_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.acc_stream_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.acc_stream_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_8_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_8_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_8_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.acc_stream_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_9_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_9_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_9_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.acc_stream_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_10_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_10_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_10_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.acc_stream_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_11_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_11_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_11_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.acc_stream_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_12_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_12_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_12_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.acc_stream_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_13_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_13_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_13_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.acc_stream_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_14_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_14_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_14_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.acc_stream_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_15_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_15_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_15_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.acc_stream_16_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_16_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_16_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_16_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.acc_stream_17_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.acc_stream_18_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.acc_stream_19_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.acc_stream_20_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.acc_stream_21_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.acc_stream_22_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.acc_stream_23_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.acc_stream_24_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    19: begin
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.start_for_conv_mukbM_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.ap_idle))) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.start_for_conv_mukbM_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_mul_U3_3.ap_idle))) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    21: begin
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.start_for_conv_aclbW_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.ap_done)) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.start_for_conv_aclbW_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.ap_done)) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    endcase
                end
                21 : begin
                    case(index2)
                    8: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.acc_stream_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.acc_stream_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.acc_stream_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.acc_stream_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.acc_stream_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.acc_stream_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.acc_stream_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.acc_stream_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.acc_stream_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_8_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_8_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_8_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.acc_stream_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_9_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_9_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_9_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.acc_stream_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_10_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_10_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_10_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.acc_stream_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_11_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_11_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_11_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.acc_stream_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_12_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_12_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_12_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.acc_stream_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_13_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_13_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_13_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.acc_stream_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_14_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_14_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_14_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.acc_stream_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_15_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_15_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_15_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.acc_stream_16_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_16_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_16_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_16_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.acc_stream_17_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.acc_stream_18_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.acc_stream_19_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.acc_stream_20_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.acc_stream_21_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.acc_stream_22_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.acc_stream_23_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.acc_stream_24_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv195_U0.grp_conv_fu_126.acc_stream_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    20: begin
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.start_for_conv_aclbW_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.ap_idle))) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.start_for_conv_aclbW_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_conv198_U0.grp_conv364_fu_126.conv_acc_U3_3.ap_idle))) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    endcase
                end
                22 : begin
                    case(index2)
                    6: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_glue_U0.grp_glue_fu_30.in_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.conv_out_0_0_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.conv_out_0_0_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.conv_out_0_0_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_vdy_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_glue_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_glue_U0.ap_idle))) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_vdy_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_glue_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_glue_U0.ap_idle))) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    10: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_glue_U0.grp_glue_fu_30.in_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.conv_out_0_1_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.conv_out_0_1_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.conv_out_0_1_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    14: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_glue_U0.grp_glue_fu_30.in_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.conv_out_0_2_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.conv_out_0_2_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.conv_out_0_2_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    18: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_glue_U0.grp_glue_fu_30.in_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.conv_out_0_3_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.conv_out_0_3_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.conv_out_0_3_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    23: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_glue_U0.grp_glue_fu_30.out_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.glue_out_0_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.glue_out_0_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.glue_out_0_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_wdI_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias199_U0.ap_done)) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_wdI_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias199_U0.ap_done)) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    24: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_glue_U0.grp_glue_fu_30.out_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.glue_out_1_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.glue_out_1_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.glue_out_1_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_xdS_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias200_U0.ap_done)) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_xdS_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias200_U0.ap_done)) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    25: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_glue_U0.grp_glue_fu_30.out_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.glue_out_2_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.glue_out_2_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.glue_out_2_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_yd2_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias201_U0.ap_done)) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_yd2_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias201_U0.ap_done)) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    26: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_glue_U0.grp_glue_fu_30.out_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.glue_out_3_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.glue_out_3_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.glue_out_3_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_zec_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias202_U0.ap_done)) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_zec_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias202_U0.ap_done)) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    endcase
                end
                23 : begin
                    case(index2)
                    22: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias199_U0.grp_bias_fu_28.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.glue_out_0_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.glue_out_0_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.glue_out_0_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_wdI_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias199_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias199_U0.ap_idle))) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_wdI_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias199_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias199_U0.ap_idle))) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    28: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias199_U0.grp_bias_fu_28.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                24 : begin
                    case(index2)
                    22: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias200_U0.grp_bias372_fu_28.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.glue_out_1_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.glue_out_1_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.glue_out_1_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_xdS_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias200_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias200_U0.ap_idle))) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_xdS_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias200_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias200_U0.ap_idle))) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    28: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias200_U0.grp_bias372_fu_28.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                25 : begin
                    case(index2)
                    22: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias201_U0.grp_bias371_fu_28.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.glue_out_2_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.glue_out_2_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.glue_out_2_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_yd2_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias201_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias201_U0.ap_idle))) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_yd2_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias201_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias201_U0.ap_idle))) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    28: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias201_U0.grp_bias371_fu_28.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                26 : begin
                    case(index2)
                    22: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias202_U0.grp_bias370_fu_28.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.glue_out_3_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.glue_out_3_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.glue_out_3_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_zec_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias202_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias202_U0.ap_idle))) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.start_for_Conv_0_zec_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias202_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias202_U0.ap_idle))) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    28: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_U0.Conv_0_bias202_U0.grp_bias370_fu_28.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                27 : begin
                    case(index2)
                    23: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_in_U0.in_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    24: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_in_U0.in_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    25: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_in_U0.in_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    26: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_in_U0.in_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    31: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    32: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    33: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    34: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    35: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    36: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    37: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    38: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    39: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_25_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_25_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_25_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    40: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_26_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_26_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_26_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    41: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_27_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_27_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_27_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    42: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_28_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_28_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_28_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    43: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_29_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_29_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_29_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    44: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_30_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_30_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_30_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    45: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_31_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_31_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_31_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    46: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_32_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_32_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_32_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    1: begin
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.start_for_Conv_0_Gfk_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.ap_idle))) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.start_for_Conv_0_Gfk_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.ap_idle))) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    30: begin
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.start_for_Relu_1_U0_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.ap_done)) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.start_for_Relu_1_U0_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.ap_done)) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    endcase
                end
                28 : begin
                    case(index2)
                    23: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_in_U0.in_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    24: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_in_U0.in_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    25: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_in_U0.in_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    26: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_in_U0.in_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_Conv_0_squeez_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    29: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_in_U0.out_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_in_U0.out_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_in_U0.out_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_in_U0.out_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_in_U0.out_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_in_U0.out_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_in_U0.out_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_in_U0.out_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_in_U0.out_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_8_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_8_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_8_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_in_U0.out_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_9_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_9_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_9_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_in_U0.out_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_10_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_10_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_10_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_in_U0.out_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_11_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_11_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_11_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_in_U0.out_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_12_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_12_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_12_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_in_U0.out_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_13_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_13_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_13_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_in_U0.out_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_14_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_14_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_14_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_in_U0.out_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_15_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_15_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_15_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.start_for_squeezeAem_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.ap_done)) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.start_for_squeezeAem_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.ap_done)) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    endcase
                end
                29 : begin
                    case(index2)
                    28: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.in_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.in_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.in_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.in_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.in_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.in_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.in_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.in_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.in_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_8_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_8_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_8_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.in_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_9_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_9_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_9_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.in_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_10_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_10_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_10_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.in_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_11_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_11_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_11_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.in_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_12_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_12_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_12_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.in_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_13_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_13_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_13_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.in_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_14_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_14_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_14_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.in_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_15_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_15_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.cache_15_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.start_for_squeezeAem_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.ap_idle))) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.start_for_squeezeAem_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.ap_idle))) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    31: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    32: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    33: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    34: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    35: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    36: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    37: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    38: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    39: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_25_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_25_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_25_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    40: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_26_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_26_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_26_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    41: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_27_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_27_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_27_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    42: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_28_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_28_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_28_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    43: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_29_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_29_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_29_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    44: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_30_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_30_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_30_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    45: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_31_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_31_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_31_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    46: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_16_U0.squeeze_U0.squeeze_out_1_U0.out_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_32_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_32_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_32_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                30 : begin
                    case(index2)
                    29: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu203_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu204_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu205_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu206_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu207_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu208_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu209_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu210_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu211_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_25_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_25_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_25_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu212_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_26_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_26_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_26_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu213_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_27_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_27_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_27_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu214_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_28_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_28_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_28_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu215_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_29_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_29_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_29_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu216_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_30_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_30_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_30_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu217_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_31_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_31_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_31_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu218_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_32_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_32_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_32_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    48: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu203_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_16_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_16_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_16_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu204_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu205_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu206_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu207_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu208_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu209_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu210_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu211_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu212_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_25_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_25_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_25_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu213_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_26_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_26_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_26_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu214_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_27_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_27_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_27_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu215_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_28_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_28_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_28_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu216_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_29_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_29_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_29_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu217_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_30_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_30_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_30_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu218_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_31_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_31_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_31_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    27: begin
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.start_for_Relu_1_U0_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.ap_idle))) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.start_for_Relu_1_U0_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.ap_idle))) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    47: begin
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.start_for_squeezeHfu_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.ap_done)) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.start_for_squeezeHfu_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.ap_done)) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    endcase
                end
                31 : begin
                    case(index2)
                    29: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu203_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    48: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu203_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_16_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_16_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_16_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                32 : begin
                    case(index2)
                    29: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu204_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    48: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu204_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                33 : begin
                    case(index2)
                    29: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu205_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    48: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu205_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                34 : begin
                    case(index2)
                    29: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu206_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    48: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu206_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                35 : begin
                    case(index2)
                    29: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu207_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    48: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu207_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                36 : begin
                    case(index2)
                    29: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu208_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    48: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu208_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                37 : begin
                    case(index2)
                    29: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu209_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    48: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu209_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                38 : begin
                    case(index2)
                    29: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu210_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    48: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu210_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                39 : begin
                    case(index2)
                    29: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu211_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_25_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_25_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_25_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    48: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu211_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                40 : begin
                    case(index2)
                    29: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu212_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_26_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_26_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_26_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    48: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu212_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_25_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_25_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_25_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                41 : begin
                    case(index2)
                    29: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu213_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_27_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_27_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_27_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    48: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu213_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_26_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_26_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_26_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                42 : begin
                    case(index2)
                    29: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu214_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_28_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_28_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_28_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    48: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu214_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_27_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_27_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_27_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                43 : begin
                    case(index2)
                    29: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu215_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_29_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_29_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_29_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    48: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu215_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_28_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_28_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_28_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                44 : begin
                    case(index2)
                    29: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu216_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_30_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_30_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_30_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    48: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu216_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_29_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_29_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_29_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                45 : begin
                    case(index2)
                    29: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu217_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_31_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_31_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_31_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    48: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu217_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_30_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_30_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_30_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                46 : begin
                    case(index2)
                    29: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu218_U0.grp_relu_fu_18.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_32_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_32_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Conv_0_squeeze_Relu_32_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    48: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_U0.Relu_1_relu218_U0.grp_relu_fu_18.out_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_31_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_31_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_31_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                47 : begin
                    case(index2)
                    31: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_16_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_16_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_16_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    32: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    33: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    34: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    35: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    36: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    37: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    38: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    39: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    40: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_25_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_25_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_25_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    41: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_26_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_26_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_26_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    42: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_27_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_27_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_27_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    43: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_28_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_28_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_28_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    44: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_29_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_29_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_29_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    45: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_30_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_30_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_30_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    46: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_31_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_31_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_31_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    50: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.out_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_0_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_0_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_0_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.out_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_1_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_1_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_1_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.out_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_2_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_2_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_2_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.out_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_3_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_3_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_3_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    30: begin
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.start_for_squeezeHfu_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.ap_idle))) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.start_for_squeezeHfu_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.ap_idle))) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    endcase
                end
                48 : begin
                    case(index2)
                    31: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_16_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_16_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_16_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    32: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_17_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_17_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_17_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    33: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_18_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_18_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_18_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    34: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_19_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_19_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_19_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    35: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_20_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_20_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_20_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    36: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_21_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_21_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_21_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    37: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_22_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_22_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_22_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    38: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_23_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_23_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_23_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    39: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_24_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_24_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_24_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    40: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_25_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_25_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_25_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    41: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_26_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_26_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_26_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    42: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_27_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_27_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_27_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    43: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_28_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_28_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_28_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    44: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_29_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_29_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_29_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    45: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_30_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_30_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_30_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    46: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.in_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_31_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_31_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.Relu_1_squeeze_Relu_31_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    49: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.out_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.out_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.out_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.out_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.out_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.out_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.out_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.out_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.out_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_8_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_8_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_8_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.out_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_9_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_9_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_9_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.out_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_10_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_10_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_10_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.out_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_11_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_11_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_11_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.out_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_12_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_12_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_12_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.out_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_13_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_13_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_13_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.out_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_14_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_14_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_14_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_in_1_U0.out_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_15_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_15_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_15_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.start_for_squeezeEe0_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.ap_done)) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.start_for_squeezeEe0_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.ap_done)) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    endcase
                end
                49 : begin
                    case(index2)
                    48: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.in_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_0_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_0_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_0_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.in_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_1_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_1_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_1_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.in_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_2_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_2_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_2_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.in_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.in_4_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_4_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_4_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_4_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.in_5_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_5_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_5_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_5_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.in_6_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_6_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_6_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_6_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.in_7_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_7_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_7_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_7_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.in_8_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_8_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_8_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_8_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.in_9_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_9_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_9_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_9_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.in_10_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_10_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_10_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_10_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.in_11_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_11_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_11_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_11_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.in_12_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_12_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_12_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_12_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.in_13_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_13_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_13_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_13_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.in_14_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_14_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_14_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_14_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.in_15_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_15_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_15_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.cache_15_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.start_for_squeezeEe0_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.ap_idle))) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.start_for_squeezeEe0_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.ap_idle))) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    50: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.out_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_0_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_0_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_0_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.out_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_1_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_1_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_1_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.out_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_2_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_2_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_2_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.squeeze_Relu_1_U0.squeeze_1_U0.squeeze_out_U0.out_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_3_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_3_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_3_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                50 : begin
                    case(index2)
                    0: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.mem_write_U0.weights_reloading_in_3_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.weights_reloading_in_3_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.weights_reloading_in_3_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.weights_reloading_in_3_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.mem_write_U0.out_hw_V_offset_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_hw_V_offset_c_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_hw_V_offset_c_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_hw_V_offset_c_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.start_for_mem_wriFfa_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.mem_write_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.mem_write_U0.ap_idle))) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.start_for_mem_wriFfa_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.mem_write_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.mem_write_U0.ap_idle))) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    49: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.mem_write_U0.out_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_0_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_0_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_0_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.mem_write_U0.out_1_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_1_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_1_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_1_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.mem_write_U0.out_2_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_2_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_2_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_2_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.mem_write_U0.out_3_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_3_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_3_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_process_r_fu_304.out_3_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                    end
                    endcase
                end
                51 : begin
                    case(index2)
                    52: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_reload_weights_fu_524.mem_read_U0.wr_0_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_reload_weights_fu_524.wr_0_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_reload_weights_fu_524.wr_0_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_reload_weights_fu_524.wr_0_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_reload_weights_fu_524.start_for_weightsbkb_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_reload_weights_fu_524.weights_reloading_U0.ap_done)) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_reload_weights_fu_524.start_for_weightsbkb_U.if_full_n & AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_reload_weights_fu_524.weights_reloading_U0.ap_done)) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    endcase
                end
                52 : begin
                    case(index2)
                    51: begin
                        if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_reload_weights_fu_524.weights_reloading_U0.in_V_V_blk_n) begin
                            chan_path = "fpgaconvnet_ip.Block_proc_U0.grp_reload_weights_fu_524.wr_0_V_V_U";
                            if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_reload_weights_fu_524.wr_0_V_V_U.if_empty_n) begin
                                $display("//      Channel: %0s, EMPTY", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_reload_weights_fu_524.wr_0_V_V_U.if_full_n) begin
                                $display("//      Channel: %0s, FULL", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                            else begin
                                $display("//      Channel: %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_path %0s", chan_path);
                                $fdisplay(fp, "Dependence_Channel_status NULL");
                            end
                        end
                        if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_reload_weights_fu_524.start_for_weightsbkb_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_reload_weights_fu_524.weights_reloading_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_reload_weights_fu_524.weights_reloading_U0.ap_idle))) begin
                            chan_path = "";
                            if ((~AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_reload_weights_fu_524.start_for_weightsbkb_U.if_empty_n & (AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_reload_weights_fu_524.weights_reloading_U0.ap_ready | AESL_inst_fpgaconvnet_ip.Block_proc_U0.grp_reload_weights_fu_524.weights_reloading_U0.ap_idle))) begin
                                $display("//      Deadlock detected: can be a false alarm due to leftover data,");
                                $display("//      please try cosim_design -disable_deadlock_detection");
                            end
                        end
                    end
                    endcase
                end
            endcase
        end
    endtask

    // report
    initial begin : report_deadlock
        integer cycle_id;
        integer cycle_comp_id;
        wait (reset == 1);
        cycle_id = 1;
        while (1) begin
            @ (negedge clock);
            case (CS_fsm)
                ST_DL_DETECTED: begin
                    cycle_comp_id = 2;
                    if (dl_detect_reg != dl_done_reg) begin
                        if (dl_done_reg == 'b0) begin
                            print_dl_head;
                        end
                        print_cycle_start(proc_path(origin), cycle_id);
                        cycle_id = cycle_id + 1;
                    end
                    else begin
                        print_dl_end(cycle_id - 1);
                        $finish;
                    end
                end
                ST_DL_REPORT: begin
                    if ((|(dl_in_vec)) & ~(|(dl_in_vec & origin_reg))) begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                        print_cycle_proc_comp(proc_path(dl_in_vec), cycle_comp_id);
                        cycle_comp_id = cycle_comp_id + 1;
                    end
                    else begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                    end
                end
            endcase
        end
    end
 
endmodule
